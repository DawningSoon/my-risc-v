module csr (
    // ports
);
    
endmodule