module ins_fetch (
    input wire [31:0]           pc_addr_i,
    input wire [31:0]           rom_inst_i
);
    
endmodule